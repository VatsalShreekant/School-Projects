library verilog;
use verilog.vl_types.all;
entity cpu1_vlg_vec_tst is
end cpu1_vlg_vec_tst;
